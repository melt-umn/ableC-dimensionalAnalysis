grammar edu:umn:cs:melt:exts:ableC:dimensionalAnalysis:concretesyntax;

exports edu:umn:cs:melt:exts:ableC:dimensionalAnalysis:concretesyntax:units;
exports edu:umn:cs:melt:exts:ableC:dimensionalAnalysis:concretesyntax:convertUnits;


