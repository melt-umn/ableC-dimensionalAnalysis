grammar edu:umn:cs:melt:exts:ableC:dimensionalAnalysis;

exports edu:umn:cs:melt:exts:ableC:dimensionalAnalysis:abstractsyntax;
exports edu:umn:cs:melt:exts:ableC:dimensionalAnalysis:concretesyntax;

