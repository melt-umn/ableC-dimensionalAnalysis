grammar edu:umn:cs:melt:exts:ableC:dimensionalAnalysis:src:concretesyntax;

exports edu:umn:cs:melt:exts:ableC:dimensionalAnalysis:src:concretesyntax:units;


