grammar edu:umn:cs:melt:exts:ableC:dimensionalAnalysis:src ;

exports edu:umn:cs:melt:exts:ableC:dimensionalAnalysis:src:abstractsyntax ;
exports edu:umn:cs:melt:exts:ableC:dimensionalAnalysis:src:concretesyntax ;

