grammar edu:umn:cs:melt:exts:ableC:dimensionalAnalysis ;

exports edu:umn:cs:melt:exts:ableC:dimensionalAnalysis:src ;

{- Exporting the 'src' directory allows extension users to simply
   place your extension directory in a directory in which they already
   keep language extensions.  This lets them easily use it in creating a
   new compiler without having to specify a path to your extension - it
   can be simply referenced by name.
 -}
