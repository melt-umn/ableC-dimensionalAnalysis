grammar edu:umn:cs:melt:exts:ableC:dimensionalAnalysis:modular_analyses:determinism;

import edu:umn:cs:melt:ableC:host only ablecParser;

copper_mda testTypeQualifier(ablecParser) {
  edu:umn:cs:melt:exts:ableC:dimensionalAnalysis:src:concretesyntax:units;
}

